module IP_encoder ();
  
endmodule
