module IP_encoder_tb ();

endmodule
